
package mem_pkg;

    import uvm_pkg::*;

    `include "uvm_macros.svh"

    `include "mem_sequence_item.svh"
    `include "mem_sequence.svh"
    `include "mem_sequencer.svh"
    `include "mem_driver.svh"
    `include "mem_monitor.svh"
    `include "mem_agent.svh"
    `include "mem_subscriber.svh"
    `include "mem_scoreboard.svh"
    `include "mem_env.svh"
    `include "mem_test.svh"
    
endpackage: mem_pkg
